module jinverter (
    y,
    a
);
    output y;
    input a;

    assign y = ~a;

endmodule
